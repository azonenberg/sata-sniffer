/***********************************************************************************************************************
*                                                                                                                      *
* sata-sniffer v0.1                                                                                                    *
*                                                                                                                      *
* Copyright (c) 2021-2022 Andrew D. Zonenberg and contributors                                                         *
* All rights reserved.                                                                                                 *
*                                                                                                                      *
* Redistribution and use in source and binary forms, with or without modification, are permitted provided that the     *
* following conditions are met:                                                                                        *
*                                                                                                                      *
*    * Redistributions of source code must retain the above copyright notice, this list of conditions, and the         *
*      following disclaimer.                                                                                           *
*                                                                                                                      *
*    * Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the       *
*      following disclaimer in the documentation and/or other materials provided with the distribution.                *
*                                                                                                                      *
*    * Neither the name of the author nor the names of any contributors may be used to endorse or promote products     *
*      derived from this software without specific prior written permission.                                           *
*                                                                                                                      *
* THIS SOFTWARE IS PROVIDED BY THE AUTHORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   *
* TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL *
* THE AUTHORS BE HELD LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES        *
* (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR       *
* BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT *
* (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE       *
* POSSIBILITY OF SUCH DAMAGE.                                                                                          *
*                                                                                                                      *
***********************************************************************************************************************/

`include "LogicPod.svh"

/**
	@brief Logic analyzer pod datapath

	This module takes in the combinatorial LVDS output of a single 8-bit logic analyzer pod (MEAD, CONWAY, etc) and
	samples it at 5 Gsps.

	All clocks must come from the same PLL and be aligned.
 */
module LogicPodDatapath #(
	parameter LANE_INVERT 	= 8'b00000000,
	parameter POD_NUMBER 	= 0
) (

	//Main clock
	input wire				clk_312p5mhz,

	//Reference clock for IDELAYs
	input wire				clk_400mhz,

	//Oversampling clocks
	input wire				clk_625mhz_fabric,
	input wire				clk_625mhz_io_0,
	input wire				clk_625mhz_io_90,

	//LVDS input
	input wire[7:0]			pod_data_p,
	input wire[7:0]			pod_data_n,

	//DDR interface
	input wire				clk_ram,
	input wire				ram_ready,
	output logic			ram_wr_en	= 0,
	output logic[28:0]		ram_wr_addr	= 0,
	output logic[255:0]		ram_wr_data	= 0,
	input wire				ram_wr_done
);

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Remap pod data lines to match front panel ordering

	wire[7:0]	pod_data_p_remapped;
	wire[7:0]	pod_data_n_remapped;

	assign pod_data_p_remapped[0] = pod_data_p[3];
	assign pod_data_n_remapped[0] = pod_data_n[3];

	assign pod_data_p_remapped[1] = pod_data_p[2];
	assign pod_data_n_remapped[1] = pod_data_n[2];

	assign pod_data_p_remapped[2] = pod_data_p[7];
	assign pod_data_n_remapped[2] = pod_data_n[7];

	assign pod_data_p_remapped[3] = pod_data_p[6];
	assign pod_data_n_remapped[3] = pod_data_n[6];

	assign pod_data_p_remapped[4] = pod_data_p[5];
	assign pod_data_n_remapped[4] = pod_data_n[5];

	assign pod_data_p_remapped[5] = pod_data_p[4];
	assign pod_data_n_remapped[5] = pod_data_n[4];

	assign pod_data_p_remapped[6] = pod_data_p[1];
	assign pod_data_n_remapped[6] = pod_data_n[1];

	assign pod_data_p_remapped[7] = pod_data_p[0];
	assign pod_data_n_remapped[7] = pod_data_n[0];

	localparam LANE_INVERT_REMAPPED =
	{
		LANE_INVERT[0],
		LANE_INVERT[1],
		LANE_INVERT[4],
		LANE_INVERT[5],
		LANE_INVERT[6],
		LANE_INVERT[7],
		LANE_INVERT[2],
		LANE_INVERT[3]
	};

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// LVDS input buffers

	wire[7:0]	data_p;
	wire[7:0]	data_n;

	for(genvar g=0; g<8; g=g+1) begin

		IBUFDS_DIFF_OUT #(
			.DIFF_TERM("TRUE"),
			.IBUF_LOW_PWR("FALSE"),
			.IOSTANDARD("LVDS")
		) ibuf (
			.I(pod_data_p_remapped[g]),
			.IB(pod_data_n_remapped[g]),
			.O(data_p[g]),
			.OB(data_n[g])
		);

	end

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Delay line calibration

	IODelayCalibration cal(.refclk(clk_400mhz));

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Input delay lines

	wire[7:0] data_p_delayed;
	wire[7:0] data_n_delayed;

	IODelayBlock #(
		.WIDTH(8),
		.CAL_FREQ(400),
		.INPUT_DELAY(00),
		.DIRECTION("IN"),
		.IS_CLOCK(0)
	) idelay_p (
		.i_pad(data_p),
		.i_fabric(data_p_delayed),

		.o_pad(),
		.o_fabric(),

		.input_en(1'b1)
	);

	IODelayBlock #(
		.WIDTH(8),
		.CAL_FREQ(400),
		.INPUT_DELAY(200),
		.DIRECTION("IN"),
		.IS_CLOCK(0)
	) idelay_n (
		.i_pad(data_n),
		.i_fabric(data_n_delayed),

		.o_pad(),
		.o_fabric(),

		.input_en(1'b1)
	);

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Initial oversampling: 4 phases of 625 MHz = 2.5 Gsps, times P and N = 5 Gsps

	wire[3:0] deser_p[7:0];
	wire[3:0] deser_n[7:0];

	logic	iserdes_rst = 0;

	//Sampling order is Q1 Q3 Q2 Q4 in oversampling mode
	//then we interleave with negative before positive
	for(genvar g=0; g<8; g=g+1) begin
		ISERDESE2 #(
			.DATA_RATE("DDR"),
			.DATA_WIDTH("4"),
			.DYN_CLKDIV_INV_EN("FALSE"),
			.DYN_CLK_INV_EN("FALSE"),
			.INTERFACE_TYPE("OVERSAMPLE"),
			.NUM_CE(1),
			.OFB_USED("FALSE"),
			.SERDES_MODE("MASTER"),
			.IOBDELAY("BOTH")
		) iserdes_p (
			.Q1(deser_p[g][0]),
			.Q2(deser_p[g][2]),
			.Q3(deser_p[g][1]),
			.Q4(deser_p[g][3]),
			.Q5(),
			.Q6(),
			.Q7(),
			.Q8(),
			.O(),
			.SHIFTOUT1(),
			.SHIFTOUT2(),
			.D(),
			.DDLY(data_p_delayed[g]),
			.CLK(clk_625mhz_io_0),
			.CLKB(!clk_625mhz_io_0),
			.CE1(1'b1),
			.CE2(1'b1),
			.RST(iserdes_rst),
			.CLKDIV(),
			.CLKDIVP(1'b0),
			.OCLK(clk_625mhz_io_90),
			.OCLKB(!clk_625mhz_io_90),
			.BITSLIP(1'b0),
			.SHIFTIN1(),
			.SHIFTIN2(),
			.OFB(),
			.DYNCLKDIVSEL(),
			.DYNCLKSEL()
		);

		ISERDESE2 #(
			.DATA_RATE("DDR"),
			.DATA_WIDTH("4"),
			.DYN_CLKDIV_INV_EN("FALSE"),
			.DYN_CLK_INV_EN("FALSE"),
			.INTERFACE_TYPE("OVERSAMPLE"),
			.NUM_CE(1),
			.OFB_USED("FALSE"),
			.SERDES_MODE("MASTER"),
			.IOBDELAY("BOTH")
		) iserdes_n (
			.Q1(deser_n[g][0]),
			.Q2(deser_n[g][2]),
			.Q3(deser_n[g][1]),
			.Q4(deser_n[g][3]),
			.Q5(),
			.Q6(),
			.Q7(),
			.Q8(),
			.O(),
			.SHIFTOUT1(),
			.SHIFTOUT2(),
			.D(),
			.DDLY(data_n_delayed[g]),
			.CLK(clk_625mhz_io_0),
			.CLKB(!clk_625mhz_io_0),
			.CE1(1'b1),
			.CE2(1'b1),
			.RST(iserdes_rst),
			.CLKDIV(),
			.CLKDIVP(1'b0),
			.OCLK(clk_625mhz_io_90),
			.OCLKB(!clk_625mhz_io_90),
			.BITSLIP(1'b0),
			.SHIFTIN1(),
			.SHIFTIN2(),
			.OFB(),
			.DYNCLKDIVSEL(),
			.DYNCLKSEL()
		);

	end

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Capturing and processing

	logic[7:0]		compressed_block_valid	= 0;
	logic[7:0]		compressed_block_clear	= 0;
	logic[254:0]	compressed_block[7:0];
	wire[10:0]		fifo_rd_size[7:0];

	for(genvar g=0; g<8; g=g+1) begin

		////////////////////////////////////////////////////////////////////////////////////////////////////////////////
		// Capture into the slow clock domain

		wire[7:0]	p_merged;
		wire[7:0]	n_merged;

		LogicPodSampling sampler (
			.clk_625mhz_fabric(clk_625mhz_fabric),
			.clk_312p5mhz(clk_312p5mhz),
			.deser_p(deser_p[g]),
			.deser_n(deser_n[g]),
			.p_out(p_merged),
			.n_out(n_merged)
		);

		////////////////////////////////////////////////////////////////////////////////////////////////////////////////
		// Merge P/N into a single 16-bit stream, inverting as necessary

		//Parallel digitized output
		la_sample_t		samples;

		//N has a larger delay than P, so it's logically earlier in the stream
		always_ff @(posedge clk_312p5mhz) begin
			for(integer i=0; i<8; i=i+1) begin
				samples.bits[i*2 + 1]	<= !n_merged[i] ^ LANE_INVERT_REMAPPED[g];
				samples.bits[i*2]		<= p_merged[i] ^ LANE_INVERT_REMAPPED[g];
			end
		end

		////////////////////////////////////////////////////////////////////////////////////////////////////////////////
		// RLE compression

		wire		compress_out_valid;
		wire		compress_out_format;
		wire[15:0]	compress_out_data;

		LogicPodCompression compressor(
			.clk(clk_312p5mhz),
			.din(samples.bits),

			.out_valid(compress_out_valid),
			.out_format(compress_out_format),
			.out_data(compress_out_data)
		);

		////////////////////////////////////////////////////////////////////////////////////////////////////////////////
		// CDC FIFO from compressor to RAM clock domain

		logic		fifo_rd_en;
		wire		fifo_rd_empty;

		logic[50:0]	fifo_wr_data	= 0;
		logic		fifo_wr_en		= 0;
		logic[1:0]	fifo_wr_phase	= 0;

		always_ff @(posedge clk_312p5mhz) begin

			fifo_wr_en					<= 0;

			//TODO: gate until memory is up
			if(compress_out_valid) begin

				fifo_wr_phase 			<= fifo_wr_phase + 1;
				if(fifo_wr_phase == 2)
					fifo_wr_phase		<= 0;

				case(fifo_wr_phase)
					0:	fifo_wr_data[50:34]	<= {compress_out_format, compress_out_data};
					1:	fifo_wr_data[33:17]	<= {compress_out_format, compress_out_data};
					default: begin
						fifo_wr_en			<= 1;
						fifo_wr_data[16:0]	<= {compress_out_format, compress_out_data};
					end
				endcase

			end

		end

		//Two block RAMs
		wire[50:0]	fifo_rd_data;
		CrossClockFifo #(
			.WIDTH(51),
			.DEPTH(1024),
			.USE_BLOCK(1),
			.OUT_REG(1)
		) cdc_fifo (

			//Write side: push in at full rate.
			//No flow control really possible here as the data can't be slowed down.
			//The FIFO will just start dropping samples if you push too fast.
			//TODO: add error flag to detect when this happens
			.wr_clk(clk_312p5mhz),
			.wr_en(fifo_wr_en),
			.wr_data(fifo_wr_data),
			.wr_size(),
			.wr_full(),
			.wr_overflow(),
			.wr_reset(1'b0),

			//Read side
			.rd_clk(clk_ram),
			.rd_en(fifo_rd_en),
			.rd_data(fifo_rd_data),
			.rd_size(fifo_rd_size[g]),
			.rd_empty(fifo_rd_empty),
			.rd_underflow(),
			.rd_reset(1'b0)
		);

		////////////////////////////////////////////////////////////////////////////////////////////////////////////////
		// Deserialization

		logic[2:0]	block_word_count	= 0;
		logic		fifo_rd_valid		= 0;

		//Pop the FIFO if we have space for it
		logic[3:0]	block_word_count_fwd;
		always_comb begin

			//Number of 51-bit words that will be valid in the buffer at the end of this cycle
			block_word_count_fwd = block_word_count + fifo_rd_valid;

			//Space in the buffer?
			fifo_rd_en	 = 0;
			if(!fifo_rd_empty) begin

				//Read if continuing an existing block, but output buffer isn't full
				if(!compressed_block_valid[g] && (block_word_count_fwd < 5))
					fifo_rd_en = 1;

				//Read if this block is done
				if(compressed_block_clear[g])
					fifo_rd_en = 1;

			end

		end

		//Data comes out of the FIFO in 34-bit words containing two compression blocks.
		//We group them 7 at a time into 238-bit blocks.
		//TODO: handle flush after we trigger (might have partial words to truncate, and partial blocks)
		always_ff @(posedge clk_ram) begin

			fifo_rd_valid					<= fifo_rd_en;
			block_word_count				<= block_word_count_fwd;

			//Handle incoming read data
			//For some reason [block_word_count] doesn't synthesize so we have to do this ugliness.
			//It still compiles to address matching and clock enables.
			if(fifo_rd_valid) begin
				for(integer i=0; i<5; i=i+1) begin
					if(block_word_count == i)
						compressed_block[g][i*51 +: 51]	<= fifo_rd_data;
				end
			end

			//Block is valid once filled
			if(block_word_count_fwd == 5)
				compressed_block_valid[g]	<= 1;

			//Block is no longer valid once consumed
			if(compressed_block_clear[g]) begin
				compressed_block_valid[g]	<= 0;
				block_word_count			<= 0;
			end

		end

	end

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Arbitration for compressed blocks into DRAM

	logic		write_valid		= 0;
	logic[2:0]	write_channel	= 0;

	wire[7:0]	block_ready		= compressed_block_valid & ~compressed_block_clear;

	always_ff @(posedge clk_ram) begin

		//Pass 1: read from highest numbered channel that's more than half full
		write_valid	= 0;
		for(integer i=0; i<8; i=i+1) begin
			if( (fifo_rd_size[i] > 512) && block_ready[i] ) begin
				write_valid	= 1;
				write_channel = i;
			end
		end

		//Pass 2: read from highest numbered channel with any data
		if(!write_valid) begin
			for(integer i=0; i<8; i=i+1) begin
				if(block_ready[i]) begin
					write_valid	= 1;
					write_channel = i;
				end
			end
		end

	end

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Main mux path

	//Each LA channel has 0x200000 (2^22) 256-bit storage locations
	logic[21:0] dram_wr_ptr[7:0];
	initial begin
		for(integer i=0; i<8; i=i+1)
			dram_wr_ptr[i] <= 0;
	end

	logic	ram_write_pending	= 0;
	always_ff @(posedge clk_ram) begin

		//Default to not writing
		ram_wr_en				<= 0;
		compressed_block_clear	<= 0;

		if(ram_wr_done)
			ram_write_pending	<= 0;

		//Something won arbitration
		if(write_valid && (!ram_write_pending || ram_wr_done)) begin
			ram_wr_en			<= 1;
			ram_write_pending	<= 1;
			ram_wr_addr			<=
			{
				1'b1,
				POD_NUMBER[0],
				write_channel,
				dram_wr_ptr[write_channel],
				2'b0
			};
			ram_wr_data			<= compressed_block[write_channel];

			dram_wr_ptr[write_channel]				<= dram_wr_ptr[write_channel] + 1;
			compressed_block_clear[write_channel]	<= 1;
		end

	end

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Debug ILA (mostly so things don't get optimized out)

	if(POD_NUMBER == 0) begin
		ila_0 ila(
			.clk(clk_ram),
			.probe0(ram_wr_en),
			.probe1(ram_wr_addr),
			.probe2(ram_wr_data),
			.probe3(compressed_block_valid),
			.probe4(compressed_block_clear),
			.probe5(fifo_rd_size[0]),
			.probe6(fifo_rd_size[1]),
			.probe7(fifo_rd_size[2]),
			.probe8(fifo_rd_size[3]),
			.probe9(fifo_rd_size[4]),
			.probe10(fifo_rd_size[5]),
			.probe11(fifo_rd_size[6]),
			.probe12(fifo_rd_size[7]),
			.probe13(write_valid),
			.probe14(write_channel),
			.probe15(block_ready),
			.probe16(ram_write_pending)
		);
	end

endmodule
